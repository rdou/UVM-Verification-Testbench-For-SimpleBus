// --------------------------------------------------------------------------------
//  SimpleBus_Vir_Base_Sequence// --------------------------------------------------------------------------------class SimpleBus_Base_Vseq extends uvm_sequence #(uvm_sequence_item);    `uvm_object_utils(SimpleBus_Base_Vseq)    SimpleBus_Bus_Sequencer #(SimpleBus_Bus_Transaction) bus_sqr_h;    SimpleBus_Dut_Sequencer #(SimpleBus_Dut_Transaction) dut_sqr_h;    function new(string name = "base_vseq");        super.new(name);    endfunctionendclass : SimpleBus_Base_Vseq// --------------------------------------------------------------------------------//  SimpleBus_Bus_Dut_Vseq// --------------------------------------------------------------------------------class SimpleBus_Bus_Dut_Vseq extends SimpleBus_Base_Vseq;    `uvm_object_utils(SimpleBus_Bus_Dut_Vseq)    SimpleBus_reg_seq bus_reg_seq;    SimpleBus_Dut_Sequence dut_seq;    function new(string name = "bus_dut_vseq");        super.new(name);    endfunction    task body();        bus_reg_seq = SimpleBus_reg_seq::type_id::create("bus_reg_seq");        dut_seq     = SimpleBus_Dut_Sequence::type_id::create("dut_seq");        fork            bus_reg_seq.start(bus_sqr_h);            dut_seq.start(dut_sqr_h);        join    endtaskendclass : SimpleBus_Bus_Dut_Vseq