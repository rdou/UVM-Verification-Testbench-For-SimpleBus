// --------------------------------------------------------------------------------
//  SimpleBus_reg_predictor
// --------------------------------------------------------------------------------
typedef uvm_reg_predictor #(SimpleBus_Bus_Transaction) SimpleBus_reg_predictor;
